// Sample Verilog Design
module design(input a, b, output y);
    assign y = a & b;
endmodule

